module ex10_top();



endmodule